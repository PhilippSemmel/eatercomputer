----------------------------------------------------------------------
-- Project      :   Eater Computer
-- Module       :   eater_top_level
-- Description  :   top level file of the eater computer
--
-- Authors      :   Philipp Semmel
-- Created      :   04.03.2023
-- Last update  :   04.03.2023
----------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY eater_top_level IS
END ENTITY eater_top_level;

ARCHITECTURE RTL OF eater_top_level IS

BEGIN
    
END ARCHITECTURE RTL;